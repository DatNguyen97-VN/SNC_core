//-----------------------------------------------
//Parameters are used to set the property of FIFO

// Default Programmable Flag Offsets
// full offset
const logic [09:00] m1 = 7;
const logic [09:00] m2 = 15;
const logic [09:00] m3 = 31;
const logic [09:00] m4 = 63;
const logic [09:00] m5 = 127;
const logic [09:00] m6 = 255;
const logic [09:00] m7 = 511;
const logic [09:00] m8 = 1023;
// empty offset
const logic [09:00] n1 = 7;
const logic [09:00] n2 = 15;
const logic [09:00] n3 = 31;
const logic [09:00] n4 = 63;
const logic [09:00] n5 = 127;
const logic [09:00] n6 = 255;
const logic [09:00] n7 = 511;
const logic [09:00] n8 = 1023;
